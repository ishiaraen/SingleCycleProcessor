module alu_tb();
		logic clk, zero;
		logic [63:0] a, b, result;
		logic [3:0] ALUControl;

		
		